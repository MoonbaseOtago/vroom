module dtbrom(input [8:0]addr, output [63:0]data);
	reg [63:0]rdata;assign data=rdata;
	always @(*)
	case (addr) // synthesis full_case parallel_case
	9'h0: rdata = 64'h79070000edfe0dd0;
	9'h1: rdata = 64'hd005000038000000;
	9'h2: rdata = 64'h1100000028000000;
	9'h3: rdata = 64'h0000000010000000;
	9'h4: rdata = 64'h98050000a9010000;
	9'h5: rdata = 64'h0000000000000000;
	9'h6: rdata = 64'h0000000000000000;
	9'h7: rdata = 64'h0000000001000000;
	9'h8: rdata = 64'h0400000003000000;
	9'h9: rdata = 64'h0200000000000000;
	9'ha: rdata = 64'h0400000003000000;
	9'hb: rdata = 64'h010000000f000000;
	9'hc: rdata = 64'h1000000003000000;
	9'hd: rdata = 64'h6e6f6f4d1b000000;
	9'he: rdata = 64'h4f52562065736142;
	9'hf: rdata = 64'h0100000000214d4f;
	9'h10: rdata = 64'h0000000073757063;
	9'h11: rdata = 64'h0400000003000000;
	9'h12: rdata = 64'h0200000000000000;
	9'h13: rdata = 64'h0400000003000000;
	9'h14: rdata = 64'h010000000f000000;
	9'h15: rdata = 64'h4075706301000000;
	9'h16: rdata = 64'h0300000000000030;
	9'h17: rdata = 64'h2100000004000000;
	9'h18: rdata = 64'h0300000000757063;
	9'h19: rdata = 64'h2d0000000c000000;
	9'h1a: rdata = 64'h0000000000000000;
	9'h1b: rdata = 64'h0300000000000000;
	9'h1c: rdata = 64'h3100000005000000;
	9'h1d: rdata = 64'h0000000079616b6f;
	9'h1e: rdata = 64'h0600000003000000;
	9'h1f: rdata = 64'h6373697238000000;
	9'h20: rdata = 64'h0300000000000076;
	9'h21: rdata = 64'h4300000009000000;
	9'h22: rdata = 64'h63616d6934367672;
	9'h23: rdata = 64'h0300000000000000;
	9'h24: rdata = 64'h4d0000000b000000;
	9'h25: rdata = 64'h76732c7663736972;
	9'h26: rdata = 64'h0300000000003933;
	9'h27: rdata = 64'h5600000004000000;
	9'h28: rdata = 64'h0300000040000000;
	9'h29: rdata = 64'h6900000004000000;
	9'h2a: rdata = 64'h0300000020000000;
	9'h2b: rdata = 64'h7600000004000000;
	9'h2c: rdata = 64'h0300000000800000;
	9'h2d: rdata = 64'h8300000004000000;
	9'h2e: rdata = 64'h0300000020000000;
	9'h2f: rdata = 64'h8e00000004000000;
	9'h30: rdata = 64'h0300000020000000;
	9'h31: rdata = 64'h9900000004000000;
	9'h32: rdata = 64'h0300000040000000;
	9'h33: rdata = 64'hac00000004000000;
	9'h34: rdata = 64'h0300000020000000;
	9'h35: rdata = 64'hb900000004000000;
	9'h36: rdata = 64'h0300000000800000;
	9'h37: rdata = 64'hc600000004000000;
	9'h38: rdata = 64'h0300000020000000;
	9'h39: rdata = 64'hd100000004000000;
	9'h3a: rdata = 64'h0300000020000000;
	9'h3b: rdata = 64'hdc00000004000000;
	9'h3c: rdata = 64'h0100000000e1f505;
	9'h3d: rdata = 64'h7075727265746e69;
	9'h3e: rdata = 64'h6f72746e6f632d74;
	9'h3f: rdata = 64'h0000000072656c6c;
	9'h40: rdata = 64'h0400000003000000;
	9'h41: rdata = 64'h01000000ec000000;
	9'h42: rdata = 64'h0000000003000000;
	9'h43: rdata = 64'h03000000fd000000;
	9'h44: rdata = 64'h380000000f000000;
	9'h45: rdata = 64'h70632c7663736972;
	9'h46: rdata = 64'h000063746e692d75;
	9'h47: rdata = 64'h0400000003000000;
	9'h48: rdata = 64'h0100000012010000;
	9'h49: rdata = 64'h0200000002000000;
	9'h4a: rdata = 64'h0100000002000000;
	9'h4b: rdata = 64'h304079726f6d656d;
	9'h4c: rdata = 64'h0300000000000000;
	9'h4d: rdata = 64'h2100000007000000;
	9'h4e: rdata = 64'h000079726f6d656d;
	9'h4f: rdata = 64'h0c00000003000000;
	9'h50: rdata = 64'h000000002d000000;
	9'h51: rdata = 64'h0000002000000000;
	9'h52: rdata = 64'h0000000003000000;
	9'h53: rdata = 64'h020000001a010000;
	9'h54: rdata = 64'h00006f6901000000;
	9'h55: rdata = 64'h0400000003000000;
	9'h56: rdata = 64'h0200000000000000;
	9'h57: rdata = 64'h0400000003000000;
	9'h58: rdata = 64'h010000000f000000;
	9'h59: rdata = 64'h0b00000003000000;
	9'h5a: rdata = 64'h706d697338000000;
	9'h5b: rdata = 64'h00007375622d656c;
	9'h5c: rdata = 64'h0000000003000000;
	9'h5d: rdata = 64'h0100000028010000;
	9'h5e: rdata = 64'h326640746e696c63;
	9'h5f: rdata = 64'h0000303030303030;
	9'h60: rdata = 64'h0d00000003000000;
	9'h61: rdata = 64'h6373697238000000;
	9'h62: rdata = 64'h30746e696c632c76;
	9'h63: rdata = 64'h0300000000000000;
	9'h64: rdata = 64'h2f01000010000000;
	9'h65: rdata = 64'h0300000001000000;
	9'h66: rdata = 64'h0700000001000000;
	9'h67: rdata = 64'h0c00000003000000;
	9'h68: rdata = 64'hffffffff2d000000;
	9'h69: rdata = 64'h00001000000000ff;
	9'h6a: rdata = 64'h0100000002000000;
	9'h6b: rdata = 64'h7075727265746e69;
	9'h6c: rdata = 64'h6f72746e6f632d74;
	9'h6d: rdata = 64'h3034664072656c6c;
	9'h6e: rdata = 64'h0000003030303030;
	9'h6f: rdata = 64'h0400000003000000;
	9'h70: rdata = 64'h01000000ec000000;
	9'h71: rdata = 64'h0000000003000000;
	9'h72: rdata = 64'h03000000fd000000;
	9'h73: rdata = 64'h380000000c000000;
	9'h74: rdata = 64'h6c702c7663736972;
	9'h75: rdata = 64'h0300000000306369;
	9'h76: rdata = 64'h4301000004000000;
	9'h77: rdata = 64'h0300000010000000;
	9'h78: rdata = 64'h2f01000010000000;
	9'h79: rdata = 64'h0900000001000000;
	9'h7a: rdata = 64'h0b00000001000000;
	9'h7b: rdata = 64'h0c00000003000000;
	9'h7c: rdata = 64'hffffffff2d000000;
	9'h7d: rdata = 64'h00000004000000f4;
	9'h7e: rdata = 64'h0400000003000000;
	9'h7f: rdata = 64'h010000004e010000;
	9'h80: rdata = 64'h0400000003000000;
	9'h81: rdata = 64'h0200000012010000;
	9'h82: rdata = 64'h0100000002000000;
	9'h83: rdata = 64'h30406c6169726573;
	9'h84: rdata = 64'h0300000000000000;
	9'h85: rdata = 64'h3800000009000000;
	9'h86: rdata = 64'h613035353631736e;
	9'h87: rdata = 64'h0300000000000000;
	9'h88: rdata = 64'h2d0000000c000000;
	9'h89: rdata = 64'h00c0ffffffffffff;
	9'h8a: rdata = 64'h0300000040000000;
	9'h8b: rdata = 64'h5f01000004000000;
	9'h8c: rdata = 64'h0300000003000000;
	9'h8d: rdata = 64'h4e01000004000000;
	9'h8e: rdata = 64'h0300000002000000;
	9'h8f: rdata = 64'h6901000004000000;
	9'h90: rdata = 64'h0300000002000000;
	9'h91: rdata = 64'hdc00000004000000;
	9'h92: rdata = 64'h02000000808d5b00;
	9'h93: rdata = 64'h6640626d01000000;
	9'h94: rdata = 64'h0030303065666666;
	9'h95: rdata = 64'h0300000003000000;
	9'h96: rdata = 64'h0000626d38000000;
	9'h97: rdata = 64'h0c00000003000000;
	9'h98: rdata = 64'hffffffff2d000000;
	9'h99: rdata = 64'h4000000000e0ffff;
	9'h9a: rdata = 64'h0400000003000000;
	9'h9b: rdata = 64'h020000004e010000;
	9'h9c: rdata = 64'h0400000003000000;
	9'h9d: rdata = 64'h0300000069010000;
	9'h9e: rdata = 64'h0400000003000000;
	9'h9f: rdata = 64'h808d5b00dc000000;
	9'ha0: rdata = 64'h0800000003000000;
	9'ha1: rdata = 64'h62616e6531000000;
	9'ha2: rdata = 64'h020000000064656c;
	9'ha3: rdata = 64'h0100000002000000;
	9'ha4: rdata = 64'h0073657361696c61;
	9'ha5: rdata = 64'h0d00000003000000;
	9'ha6: rdata = 64'h2f6f692f74010000;
	9'ha7: rdata = 64'h30406c6169726573;
	9'ha8: rdata = 64'h0200000000000000;
	9'ha9: rdata = 64'h736f686301000000;
	9'haa: rdata = 64'h0300000000006e65;
	9'hab: rdata = 64'h7a0100000f000000;
	9'hac: rdata = 64'h31313a3074726175;
	9'had: rdata = 64'h0000386e30303235;
	9'hae: rdata = 64'h2700000003000000;
	9'haf: rdata = 64'h736e6f6386010000;
	9'hb0: rdata = 64'h537974743d656c6f;
	9'hb1: rdata = 64'h3030323531312c30;
	9'hb2: rdata = 64'h2067756265642020;
	9'hb3: rdata = 64'h6c6576656c676f6c;
	9'hb4: rdata = 64'h020000000000373d;
	9'hb5: rdata = 64'h666e6f6301000000;
	9'hb6: rdata = 64'h0300000000006769;
	9'hb7: rdata = 64'h8f01000004000000;
	9'hb8: rdata = 64'h0200000000501000;
	9'hb9: rdata = 64'h0900000002000000;
	9'hba: rdata = 64'h7373657264646123;
	9'hbb: rdata = 64'h2300736c6c65632d;
	9'hbc: rdata = 64'h6c65632d657a6973;
	9'hbd: rdata = 64'h6c65646f6d00736c;
	9'hbe: rdata = 64'h5f65636976656400;
	9'hbf: rdata = 64'h6765720065707974;
	9'hc0: rdata = 64'h0073757461747300;
	9'hc1: rdata = 64'h62697461706d6f63;
	9'hc2: rdata = 64'h766373697200656c;
	9'hc3: rdata = 64'h756d6d006173692c;
	9'hc4: rdata = 64'h2d6900657079742d;
	9'hc5: rdata = 64'h6c622d6568636163;
	9'hc6: rdata = 64'h657a69732d6b636f;
	9'hc7: rdata = 64'h65686361632d6900;
	9'hc8: rdata = 64'h2d6900737465732d;
	9'hc9: rdata = 64'h69732d6568636163;
	9'hca: rdata = 64'h626c742d6900657a;
	9'hcb: rdata = 64'h2d6900737465732d;
	9'hcc: rdata = 64'h657a69732d626c74;
	9'hcd: rdata = 64'h65686361632d6400;
	9'hce: rdata = 64'h732d6b636f6c622d;
	9'hcf: rdata = 64'h61632d6400657a69;
	9'hd0: rdata = 64'h737465732d656863;
	9'hd1: rdata = 64'h65686361632d6400;
	9'hd2: rdata = 64'h2d6400657a69732d;
	9'hd3: rdata = 64'h737465732d626c74;
	9'hd4: rdata = 64'h732d626c742d6400;
	9'hd5: rdata = 64'h636f6c6300657a69;
	9'hd6: rdata = 64'h6575716572662d6b;
	9'hd7: rdata = 64'h746e69230079636e;
	9'hd8: rdata = 64'h632d747075727265;
	9'hd9: rdata = 64'h746e6900736c6c65;
	9'hda: rdata = 64'h632d747075727265;
	9'hdb: rdata = 64'h656c6c6f72746e6f;
	9'hdc: rdata = 64'h6c646e6168700072;
	9'hdd: rdata = 64'h746f6f622d750065;
	9'hde: rdata = 64'h006c70732d6d642c;
	9'hdf: rdata = 64'h69007365676e6172;
	9'he0: rdata = 64'h747075727265746e;
	9'he1: rdata = 64'h646e657478652d73;
	9'he2: rdata = 64'h7663736972006465;
	9'he3: rdata = 64'h6e69007665646e2c;
	9'he4: rdata = 64'h2d74707572726574;
	9'he5: rdata = 64'h7200746e65726170;
	9'he6: rdata = 64'h74666968732d6765;
	9'he7: rdata = 64'h75727265746e6900;
	9'he8: rdata = 64'h7472617500737470;
	9'he9: rdata = 64'h74756f6474730030;
	9'hea: rdata = 64'h6f6200687461702d;
	9'heb: rdata = 64'h750073677261746f;
	9'hec: rdata = 64'h70732c746f6f622d;
	9'hed: rdata = 64'h616f6c7961702d6c;
	9'hee: rdata = 64'h74657366666f2d64;
	9'hef: rdata = 64'h74657366666f2d00;

	endcase
endmodule
